// Modulo de memoria de programa 
module dmem(input clk, mem_write,
				input  [31:0] addr,
				input  [16:0] vaddr,
				input  [31:0] write_data,
				output [31:0] read_data,
				output [7:0] vdata);

  reg [31:0] RAM[76799:0];

  initial
  begin
    RAM[212] = 8'b00111111; // .video
    RAM[213] = 8'b00111111;
    RAM[214] = 8'b00111111;
    RAM[215] = 8'b00111111;
    RAM[216] = 8'b00111111;
    RAM[217] = 8'b00111111;
    RAM[218] = 8'b00111111;
    RAM[219] = 8'b00110000;
    RAM[220] = 8'b00110000;
    RAM[221] = 8'b00110000;
    RAM[222] = 8'b00110000;
    RAM[223] = 8'b00110000;
    RAM[224] = 8'b00111111;
    RAM[225] = 8'b00111111;
    RAM[226] = 8'b00111000;
    RAM[227] = 8'b00111000;
    RAM[228] = 8'b00111000;
    RAM[229] = 8'b00111111;
    RAM[230] = 8'b00111111;
    RAM[231] = 8'b00111111;
    RAM[232] = 8'b00111111;
    RAM[233] = 8'b00111111;
    RAM[234] = 8'b00111111;
    RAM[235] = 8'b00111111;
    RAM[236] = 8'b00111111;
    RAM[237] = 8'b00111111;
    RAM[238] = 8'b00110000;
    RAM[239] = 8'b00110000;
    RAM[240] = 8'b00110000;
    RAM[241] = 8'b00110000;
    RAM[242] = 8'b00110000;
    RAM[243] = 8'b00110000;
    RAM[244] = 8'b00110000;
    RAM[245] = 8'b00110000;
    RAM[246] = 8'b00110000;
    RAM[247] = 8'b00111000;
    RAM[248] = 8'b00111000;
    RAM[249] = 8'b00111111;
    RAM[250] = 8'b00111111;
    RAM[251] = 8'b00111111;
    RAM[252] = 8'b00111111;
    RAM[253] = 8'b00111111;
    RAM[254] = 8'b00111111;
    RAM[255] = 8'b00111111;
    RAM[256] = 8'b00111111;
    RAM[257] = 8'b00111111;
    RAM[258] = 8'b00010000;
    RAM[259] = 8'b00010000;
    RAM[260] = 8'b00010000;
    RAM[261] = 8'b00111000;
    RAM[262] = 8'b00111000;
    RAM[263] = 8'b00000000;
    RAM[264] = 8'b00111000;
    RAM[265] = 8'b00110000;
    RAM[266] = 8'b00110000;
    RAM[267] = 8'b00110000;
    RAM[268] = 8'b00110000;
    RAM[269] = 8'b00111111;
    RAM[270] = 8'b00111111;
    RAM[271] = 8'b00111111;
    RAM[272] = 8'b00111111;
    RAM[273] = 8'b00111111;
    RAM[274] = 8'b00111111;
    RAM[275] = 8'b00111111;
    RAM[276] = 8'b00111111;
    RAM[277] = 8'b00010000;
    RAM[278] = 8'b00111000;
    RAM[279] = 8'b00010000;
    RAM[280] = 8'b00111000;
    RAM[281] = 8'b00111000;
    RAM[282] = 8'b00111000;
    RAM[283] = 8'b00000000;
    RAM[284] = 8'b00111000;
    RAM[285] = 8'b00111000;
    RAM[286] = 8'b00111000;
    RAM[287] = 8'b00110000;
    RAM[288] = 8'b00110000;
    RAM[289] = 8'b00111111;
    RAM[290] = 8'b00111111;
    RAM[291] = 8'b00111111;
    RAM[292] = 8'b00111111;
    RAM[293] = 8'b00111111;
    RAM[294] = 8'b00111111;
    RAM[295] = 8'b00111111;
    RAM[296] = 8'b00111111;
    RAM[297] = 8'b00010000;
    RAM[298] = 8'b00111000;
    RAM[299] = 8'b00010000;
    RAM[300] = 8'b00010000;
    RAM[301] = 8'b00111000;
    RAM[302] = 8'b00111000;
    RAM[303] = 8'b00111000;
    RAM[304] = 8'b00000000;
    RAM[305] = 8'b00111000;
    RAM[306] = 8'b00111000;
    RAM[307] = 8'b00111000;
    RAM[308] = 8'b00110000;
    RAM[309] = 8'b00111111;
    RAM[310] = 8'b00111111;
    RAM[311] = 8'b00111111;
    RAM[312] = 8'b00111111;
    RAM[313] = 8'b00111111;
    RAM[314] = 8'b00111111;
    RAM[315] = 8'b00111111;
    RAM[316] = 8'b00111111;
    RAM[317] = 8'b00010000;
    RAM[318] = 8'b00010000;
    RAM[319] = 8'b00111000;
    RAM[320] = 8'b00111000;
    RAM[321] = 8'b00111000;
    RAM[322] = 8'b00111000;
    RAM[323] = 8'b00000000;
    RAM[324] = 8'b00000000;
    RAM[325] = 8'b00000000;
    RAM[326] = 8'b00000000;
    RAM[327] = 8'b00000000;
    RAM[328] = 8'b00111111;
    RAM[329] = 8'b00111111;
    RAM[330] = 8'b00111111;
    RAM[331] = 8'b00111111;
    RAM[332] = 8'b00111111;
    RAM[333] = 8'b00111111;
    RAM[334] = 8'b00111111;
    RAM[335] = 8'b00111111;
    RAM[336] = 8'b00111111;
    RAM[337] = 8'b00111111;
    RAM[338] = 8'b00111111;
    RAM[339] = 8'b00111000;
    RAM[340] = 8'b00111000;
    RAM[341] = 8'b00111000;
    RAM[342] = 8'b00111000;
    RAM[343] = 8'b00111000;
    RAM[344] = 8'b00111000;
    RAM[345] = 8'b00111000;
    RAM[346] = 8'b00110000;
    RAM[347] = 8'b00110000;
    RAM[348] = 8'b00111111;
    RAM[349] = 8'b00111111;
    RAM[350] = 8'b00111111;
    RAM[351] = 8'b00111111;
    RAM[352] = 8'b00111111;
    RAM[353] = 8'b00111111;
    RAM[354] = 8'b00111111;
    RAM[355] = 8'b00111111;
    RAM[356] = 8'b00110000;
    RAM[357] = 8'b00110000;
    RAM[358] = 8'b00110000;
    RAM[359] = 8'b00110000;
    RAM[360] = 8'b00000011;
    RAM[361] = 8'b00110000;
    RAM[362] = 8'b00110000;
    RAM[363] = 8'b00110000;
    RAM[364] = 8'b00000011;
    RAM[365] = 8'b00110000;
    RAM[366] = 8'b00110000;
    RAM[367] = 8'b00111111;
    RAM[368] = 8'b00111111;
    RAM[369] = 8'b00010000;
    RAM[370] = 8'b00111111;
    RAM[371] = 8'b00111111;
    RAM[372] = 8'b00111111;
    RAM[373] = 8'b00111111;
    RAM[374] = 8'b00111000;
    RAM[375] = 8'b00111000;
    RAM[376] = 8'b00110000;
    RAM[377] = 8'b00110000;
    RAM[378] = 8'b00110000;
    RAM[379] = 8'b00110000;
    RAM[380] = 8'b00110000;
    RAM[381] = 8'b00000011;
    RAM[382] = 8'b00110000;
    RAM[383] = 8'b00110000;
    RAM[384] = 8'b00110000;
    RAM[385] = 8'b00000011;
    RAM[386] = 8'b00111111;
    RAM[387] = 8'b00111111;
    RAM[388] = 8'b00010000;
    RAM[389] = 8'b00010000;
    RAM[390] = 8'b00111111;
    RAM[391] = 8'b00111111;
    RAM[392] = 8'b00111111;
    RAM[393] = 8'b00111111;
    RAM[394] = 8'b00111000;
    RAM[395] = 8'b00111000;
    RAM[396] = 8'b00111000;
    RAM[397] = 8'b00110000;
    RAM[398] = 8'b00110000;
    RAM[399] = 8'b00110000;
    RAM[400] = 8'b00110000;
    RAM[401] = 8'b00000011;
    RAM[402] = 8'b00000011;
    RAM[403] = 8'b00000011;
    RAM[404] = 8'b00000011;
    RAM[405] = 8'b00111100;
    RAM[406] = 8'b00000011;
    RAM[407] = 8'b00000011;
    RAM[408] = 8'b00010000;
    RAM[409] = 8'b00010000;
    RAM[410] = 8'b00111111;
    RAM[411] = 8'b00111111;
    RAM[412] = 8'b00111111;
    RAM[413] = 8'b00111111;
    RAM[414] = 8'b00111111;
    RAM[415] = 8'b00111000;
    RAM[416] = 8'b00111111;
    RAM[417] = 8'b00111111;
    RAM[418] = 8'b00000011;
    RAM[419] = 8'b00000011;
    RAM[420] = 8'b00000011;
    RAM[421] = 8'b00000011;
    RAM[422] = 8'b00111100;
    RAM[423] = 8'b00000011;
    RAM[424] = 8'b00000011;
    RAM[425] = 8'b00000011;
    RAM[426] = 8'b00000011;
    RAM[427] = 8'b00000011;
    RAM[428] = 8'b00010000;
    RAM[429] = 8'b00010000;
    RAM[430] = 8'b00111111;
    RAM[431] = 8'b00111111;
    RAM[432] = 8'b00111111;
    RAM[433] = 8'b00111111;
    RAM[434] = 8'b00111111;
    RAM[435] = 8'b00111111;
    RAM[436] = 8'b00010000;
    RAM[437] = 8'b00010000;
    RAM[438] = 8'b00000011;
    RAM[439] = 8'b00000011;
    RAM[440] = 8'b00000011;
    RAM[441] = 8'b00000011;
    RAM[442] = 8'b00000011;
    RAM[443] = 8'b00000011;
    RAM[444] = 8'b00000011;
    RAM[445] = 8'b00000011;
    RAM[446] = 8'b00000011;
    RAM[447] = 8'b00000011;
    RAM[448] = 8'b00010000;
    RAM[449] = 8'b00010000;
    RAM[450] = 8'b00111111;
    RAM[451] = 8'b00111111;
    RAM[452] = 8'b00111111;
    RAM[453] = 8'b00111111;
    RAM[454] = 8'b00111111;
    RAM[455] = 8'b00010000;
    RAM[456] = 8'b00010000;
    RAM[457] = 8'b00010000;
    RAM[458] = 8'b00000011;
    RAM[459] = 8'b00000011;
    RAM[460] = 8'b00000011;
    RAM[461] = 8'b00000011;
    RAM[462] = 8'b00000011;
    RAM[463] = 8'b00000011;
    RAM[464] = 8'b00111111;
    RAM[465] = 8'b00111111;
    RAM[466] = 8'b00111111;
    RAM[467] = 8'b00111111;
    RAM[468] = 8'b00111111;
    RAM[469] = 8'b00111111;
    RAM[470] = 8'b00111111;
    RAM[471] = 8'b00111111;
    RAM[472] = 8'b00111111;
    RAM[473] = 8'b00111111;
    RAM[474] = 8'b00111111;
    RAM[475] = 8'b00010000;
    RAM[476] = 8'b00010000;
    RAM[477] = 8'b00111111;
    RAM[478] = 8'b00111111;
    RAM[479] = 8'b00111111;
    RAM[480] = 8'b00111111;
    RAM[481] = 8'b00111111;
    RAM[482] = 8'b00111111;
    RAM[483] = 8'b00111111;
    RAM[484] = 8'b00111111;
    RAM[485] = 8'b00111111;
    RAM[486] = 8'b00111111;
    RAM[487] = 8'b00111111;
    RAM[488] = 8'b00111111;
    RAM[489] = 8'b00111111;
    RAM[490] = 8'b00111111;
    RAM[491] = 8'b00111111;
    RAM[492] = 8'b00111111;
    RAM[493] = 8'b00111111;
    RAM[494] = 8'b00111111;
    RAM[495] = 8'b00111111;
    RAM[496] = 8'b00111111;
    RAM[497] = 8'b00111111;
    RAM[498] = 8'b00111111;
    RAM[499] = 8'b00111111;
    RAM[500] = 8'b00111111;
    RAM[501] = 8'b00111111;
    RAM[502] = 8'b00111111;
    RAM[503] = 8'b00111111;
    RAM[504] = 8'b00111111;
    RAM[505] = 8'b00111111;
    RAM[506] = 8'b00000011;
    RAM[507] = 8'b00001100;
    RAM[508] = 8'b00110000;
    RAM[509] = 8'b00111100;
    RAM[510] = 8'b00110011;
    RAM[511] = 8'b00001111;
  end

  assign vdata = RAM[{23'b0, vaddr}]; 
  assign read_data = RAM[addr[31:0]]; // word aligned
  
  always_ff @(posedge clk) 
    if (mem_write) 
	 begin
		RAM[addr[31:0]] <= write_data;
	end
endmodule


// Modulo de memoria das instruçoes
module imem(input  logic [31:0] pc,
            output logic [31:0] instr);

  logic [31:0] RAM[16:0];

  initial
  begin
		RAM[0 ]  = 32'h00000293;
		RAM[1 ]	= 32'h12c00313;
		RAM[2 ]	= 32'h00028023;
		RAM[3 ]	= 32'h00128293;
		RAM[4 ]	= 32'h0062d463;
		RAM[5 ]	= 32'hff5ff06f;
		RAM[6 ]	= 32'h0000006f;
  end

  assign instr = RAM[pc[31:2]]; // word aligned
endmodule