// Modulo de memoria de programa 
module dmem(input clk, mem_write,
				input  [31:0] addr, vaddr, write_data,
				output [31:0] read_data,
				output [31:0] vdata);

  reg [31:0] RAM[1000:0];

  initial
  begin
    RAM[0] =	32'b00000000000000000000000000111111;
    RAM[1] =	32'b00000000000000000000000000111111;
    RAM[2] =	32'b00000000000000000000000000111111;
    RAM[3] =	32'b00000000000000000000000000111111;
    RAM[4] =	32'b00000000000000000000000000111111;
    RAM[5] =	32'b00000000000000000000000000111111;
    RAM[6] =	32'b00000000000000000000000000111111;
    RAM[7] =	32'b00000000000000000000000000110000;
    RAM[8] =	32'b00000000000000000000000000110000;
    RAM[9] =	32'b00000000000000000000000000110000;
    RAM[10] =	32'b00000000000000000000000000110000;
    RAM[11] =	32'b00000000000000000000000000110000;
    RAM[12] =	32'b00000000000000000000000000111111;
    RAM[13] =	32'b00000000000000000000000000111111;
    RAM[14] =	32'b00000000000000000000000000111000;
    RAM[15] =	32'b00000000000000000000000000111000;
    RAM[16] =	32'b00000000000000000000000000111000;
    RAM[17] =	32'b00000000000000000000000000111111;
    RAM[18] =	32'b00000000000000000000000000111111;
    RAM[19] =	32'b00000000000000000000000000111111;
    RAM[20] =	32'b00000000000000000000000000111111;
    RAM[21] =	32'b00000000000000000000000000111111;
    RAM[22] =	32'b00000000000000000000000000111111;
    RAM[23] =	32'b00000000000000000000000000111111;
    RAM[24] =	32'b00000000000000000000000000111111;
    RAM[25] =	32'b00000000000000000000000000111111;
    RAM[26] =	32'b00000000000000000000000000110000;
    RAM[27] =	32'b00000000000000000000000000110000;
    RAM[28] =	32'b00000000000000000000000000110000;
    RAM[29] =	32'b00000000000000000000000000110000;
    RAM[30] =	32'b00000000000000000000000000110000;
    RAM[31] =	32'b00000000000000000000000000110000;
    RAM[32] =	32'b00000000000000000000000000110000;
    RAM[33] =	32'b00000000000000000000000000110000;
    RAM[34] =	32'b00000000000000000000000000110000;
    RAM[35] =	32'b00000000000000000000000000111000;
    RAM[36] =	32'b00000000000000000000000000111000;
    RAM[37] =	32'b00000000000000000000000000111111;
    RAM[38] =	32'b00000000000000000000000000111111;
    RAM[39] =	32'b00000000000000000000000000111111;
    RAM[40] =	32'b00000000000000000000000000111111;
    RAM[41] =	32'b00000000000000000000000000111111;
    RAM[42] =	32'b00000000000000000000000000111111;
    RAM[43] =	32'b00000000000000000000000000111111;
    RAM[44] =	32'b00000000000000000000000000111111;
    RAM[45] =	32'b00000000000000000000000000111111;
    RAM[46] =	32'b00000000000000000000000000010000;
    RAM[47] =	32'b00000000000000000000000000010000;
    RAM[48] =	32'b00000000000000000000000000010000;
    RAM[49] =	32'b00000000000000000000000000111000;
    RAM[50] =	32'b00000000000000000000000000111000;
    RAM[51] =	32'b00000000000000000000000000000000;
    RAM[52] =	32'b00000000000000000000000000111000;
    RAM[53] =	32'b00000000000000000000000000110000;
    RAM[54] =	32'b00000000000000000000000000110000;
    RAM[55] =	32'b00000000000000000000000000110000;
    RAM[56] =	32'b00000000000000000000000000110000;
    RAM[57] =	32'b00000000000000000000000000111111;
    RAM[58] =	32'b00000000000000000000000000111111;
    RAM[59] =	32'b00000000000000000000000000111111;
    RAM[60] =	32'b00000000000000000000000000111111;
    RAM[61] =	32'b00000000000000000000000000111111;
    RAM[62] =	32'b00000000000000000000000000111111;
    RAM[63] =	32'b00000000000000000000000000111111;
    RAM[64] =	32'b00000000000000000000000000111111;
    RAM[65] =	32'b00000000000000000000000000010000;
    RAM[66] =	32'b00000000000000000000000000111000;
    RAM[67] =	32'b00000000000000000000000000010000;
    RAM[68] =	32'b00000000000000000000000000111000;
    RAM[69] =	32'b00000000000000000000000000111000;
    RAM[70] =	32'b00000000000000000000000000111000;
    RAM[71] =	32'b00000000000000000000000000000000;
    RAM[72] =	32'b00000000000000000000000000111000;
    RAM[73] =	32'b00000000000000000000000000111000;
    RAM[74] =	32'b00000000000000000000000000111000;
    RAM[75] =	32'b00000000000000000000000000110000;
    RAM[76] =	32'b00000000000000000000000000110000;
    RAM[77] =	32'b00000000000000000000000000111111;
    RAM[78] =	32'b00000000000000000000000000111111;
    RAM[79] =	32'b00000000000000000000000000111111;
    RAM[80] =	32'b00000000000000000000000000111111;
    RAM[81] =	32'b00000000000000000000000000111111;
    RAM[82] =	32'b00000000000000000000000000111111;
    RAM[83] =	32'b00000000000000000000000000111111;
    RAM[84] =	32'b00000000000000000000000000111111;
    RAM[85] =	32'b00000000000000000000000000010000;
    RAM[86] =	32'b00000000000000000000000000111000;
    RAM[87] =	32'b00000000000000000000000000010000;
    RAM[88] =	32'b00000000000000000000000000010000;
    RAM[89] =	32'b00000000000000000000000000111000;
    RAM[90] =	32'b00000000000000000000000000111000;
    RAM[91] =	32'b00000000000000000000000000111000;
    RAM[92] =	32'b00000000000000000000000000000000;
    RAM[93] =	32'b00000000000000000000000000111000;
    RAM[94] =	32'b00000000000000000000000000111000;
    RAM[95] =	32'b00000000000000000000000000111000;
    RAM[96] =	32'b00000000000000000000000000110000;
    RAM[97] =	32'b00000000000000000000000000111111;
    RAM[98] =	32'b00000000000000000000000000111111;
    RAM[99] =	32'b00000000000000000000000000111111;
    RAM[100] =	32'b00000000000000000000000000111111;
    RAM[101] =	32'b00000000000000000000000000111111;
    RAM[102] =	32'b00000000000000000000000000111111;
    RAM[103] =	32'b00000000000000000000000000111111;
    RAM[104] =	32'b00000000000000000000000000111111;
    RAM[105] =	32'b00000000000000000000000000010000;
    RAM[106] =	32'b00000000000000000000000000010000;
    RAM[107] =	32'b00000000000000000000000000111000;
    RAM[108] =	32'b00000000000000000000000000111000;
    RAM[109] =	32'b00000000000000000000000000111000;
    RAM[110] =	32'b00000000000000000000000000111000;
    RAM[111] =	32'b00000000000000000000000000000000;
    RAM[112] =	32'b00000000000000000000000000000000;
    RAM[113] =	32'b00000000000000000000000000000000;
    RAM[114] =	32'b00000000000000000000000000000000;
    RAM[115] =	32'b00000000000000000000000000000000;
    RAM[116] =	32'b00000000000000000000000000111111;
    RAM[117] =	32'b00000000000000000000000000111111;
    RAM[118] =	32'b00000000000000000000000000111111;
    RAM[119] =	32'b00000000000000000000000000111111;
    RAM[120] =	32'b00000000000000000000000000111111;
    RAM[121] =	32'b00000000000000000000000000111111;
    RAM[122] =	32'b00000000000000000000000000111111;
    RAM[123] =	32'b00000000000000000000000000111111;
    RAM[124] =	32'b00000000000000000000000000111111;
    RAM[125] =	32'b00000000000000000000000000111111;
    RAM[126] =	32'b00000000000000000000000000111111;
    RAM[127] =	32'b00000000000000000000000000111000;
    RAM[128] =	32'b00000000000000000000000000111000;
    RAM[129] =	32'b00000000000000000000000000111000;
    RAM[130] =	32'b00000000000000000000000000111000;
    RAM[131] =	32'b00000000000000000000000000111000;
    RAM[132] =	32'b00000000000000000000000000111000;
    RAM[133] =	32'b00000000000000000000000000111000;
    RAM[134] =	32'b00000000000000000000000000110000;
    RAM[135] =	32'b00000000000000000000000000110000;
    RAM[136] =	32'b00000000000000000000000000111111;
    RAM[137] =	32'b00000000000000000000000000111111;
    RAM[138] =	32'b00000000000000000000000000111111;
    RAM[139] =	32'b00000000000000000000000000111111;
    RAM[140] =	32'b00000000000000000000000000111111;
    RAM[141] =	32'b00000000000000000000000000111111;
    RAM[142] =	32'b00000000000000000000000000111111;
    RAM[143] =	32'b00000000000000000000000000111111;
    RAM[144] =	32'b00000000000000000000000000110000;
    RAM[145] =	32'b00000000000000000000000000110000;
    RAM[146] =	32'b00000000000000000000000000110000;
    RAM[147] =	32'b00000000000000000000000000110000;
    RAM[148] =	32'b00000000000000000000000000000011;
    RAM[149] =	32'b00000000000000000000000000110000;
    RAM[150] =	32'b00000000000000000000000000110000;
    RAM[151] =	32'b00000000000000000000000000110000;
    RAM[152] =	32'b00000000000000000000000000000011;
    RAM[153] =	32'b00000000000000000000000000110000;
    RAM[154] =	32'b00000000000000000000000000110000;
    RAM[155] =	32'b00000000000000000000000000111111;
    RAM[156] =	32'b00000000000000000000000000111111;
    RAM[157] =	32'b00000000000000000000000000010000;
    RAM[158] =	32'b00000000000000000000000000111111;
    RAM[159] =	32'b00000000000000000000000000111111;
    RAM[160] =	32'b00000000000000000000000000111111;
    RAM[161] =	32'b00000000000000000000000000111111;
    RAM[162] =	32'b00000000000000000000000000111000;
    RAM[163] =	32'b00000000000000000000000000111000;
    RAM[164] =	32'b00000000000000000000000000110000;
    RAM[165] =	32'b00000000000000000000000000110000;
    RAM[166] =	32'b00000000000000000000000000110000;
    RAM[167] =	32'b00000000000000000000000000110000;
    RAM[168] =	32'b00000000000000000000000000110000;
    RAM[169] =	32'b00000000000000000000000000000011;
    RAM[170] =	32'b00000000000000000000000000110000;
    RAM[171] =	32'b00000000000000000000000000110000;
    RAM[172] =	32'b00000000000000000000000000110000;
    RAM[173] =	32'b00000000000000000000000000000011;
    RAM[174] =	32'b00000000000000000000000000111111;
    RAM[175] =	32'b00000000000000000000000000111111;
    RAM[176] =	32'b00000000000000000000000000010000;
    RAM[177] =	32'b00000000000000000000000000010000;
    RAM[178] =	32'b00000000000000000000000000111111;
    RAM[179] =	32'b00000000000000000000000000111111;
    RAM[180] =	32'b00000000000000000000000000111111;
    RAM[181] =	32'b00000000000000000000000000111111;
    RAM[182] =	32'b00000000000000000000000000111000;
    RAM[183] =	32'b00000000000000000000000000111000;
    RAM[184] =	32'b00000000000000000000000000111000;
    RAM[185] =	32'b00000000000000000000000000110000;
    RAM[186] =	32'b00000000000000000000000000110000;
    RAM[187] =	32'b00000000000000000000000000110000;
    RAM[188] =	32'b00000000000000000000000000110000;
    RAM[189] =	32'b00000000000000000000000000000011;
    RAM[190] =	32'b00000000000000000000000000000011;
    RAM[191] =	32'b00000000000000000000000000000011;
    RAM[192] =	32'b00000000000000000000000000000011;
    RAM[193] =	32'b00000000000000000000000000111100;
    RAM[194] =	32'b00000000000000000000000000000011;
    RAM[195] =	32'b00000000000000000000000000000011;
    RAM[196] =	32'b00000000000000000000000000010000;
    RAM[197] =	32'b00000000000000000000000000010000;
    RAM[198] =	32'b00000000000000000000000000111111;
    RAM[199] =	32'b00000000000000000000000000111111;
    RAM[200] =	32'b00000000000000000000000000111111;
    RAM[201] =	32'b00000000000000000000000000111111;
    RAM[202] =	32'b00000000000000000000000000111111;
    RAM[203] =	32'b00000000000000000000000000111000;
    RAM[204] =	32'b00000000000000000000000000111111;
    RAM[205] =	32'b00000000000000000000000000111111;
    RAM[206] =	32'b00000000000000000000000000000011;
    RAM[207] =	32'b00000000000000000000000000000011;
    RAM[208] =	32'b00000000000000000000000000000011;
    RAM[209] =	32'b00000000000000000000000000000011;
    RAM[210] =	32'b00000000000000000000000000111100;
    RAM[211] =	32'b00000000000000000000000000000011;
    RAM[212] =	32'b00000000000000000000000000000011;
    RAM[213] =	32'b00000000000000000000000000000011;
    RAM[214] =	32'b00000000000000000000000000000011;
    RAM[215] =	32'b00000000000000000000000000000011;
    RAM[216] =	32'b00000000000000000000000000010000;
    RAM[217] =	32'b00000000000000000000000000010000;
    RAM[218] =	32'b00000000000000000000000000111111;
    RAM[219] =	32'b00000000000000000000000000111111;
    RAM[220] =	32'b00000000000000000000000000111111;
    RAM[221] =	32'b00000000000000000000000000111111;
    RAM[222] =	32'b00000000000000000000000000111111;
    RAM[223] =	32'b00000000000000000000000000111111;
    RAM[224] =	32'b00000000000000000000000000010000;
    RAM[225] =	32'b00000000000000000000000000010000;
    RAM[226] =	32'b00000000000000000000000000000011;
    RAM[227] =	32'b00000000000000000000000000000011;
    RAM[228] =	32'b00000000000000000000000000000011;
    RAM[229] =	32'b00000000000000000000000000000011;
    RAM[230] =	32'b00000000000000000000000000000011;
    RAM[231] =	32'b00000000000000000000000000000011;
    RAM[232] =	32'b00000000000000000000000000000011;
    RAM[233] =	32'b00000000000000000000000000000011;
    RAM[234] =	32'b00000000000000000000000000000011;
    RAM[235] =	32'b00000000000000000000000000000011;
    RAM[236] =	32'b00000000000000000000000000010000;
    RAM[237] =	32'b00000000000000000000000000010000;
    RAM[238] =	32'b00000000000000000000000000111111;
    RAM[239] =	32'b00000000000000000000000000111111;
    RAM[240] =	32'b00000000000000000000000000111111;
    RAM[241] =	32'b00000000000000000000000000111111;
    RAM[242] =	32'b00000000000000000000000000111111;
    RAM[243] =	32'b00000000000000000000000000010000;
    RAM[244] =	32'b00000000000000000000000000010000;
    RAM[245] =	32'b00000000000000000000000000010000;
    RAM[246] =	32'b00000000000000000000000000000011;
    RAM[247] =	32'b00000000000000000000000000000011;
    RAM[248] =	32'b00000000000000000000000000000011;
    RAM[249] =	32'b00000000000000000000000000000011;
    RAM[250] =	32'b00000000000000000000000000000011;
    RAM[251] =	32'b00000000000000000000000000000011;
    RAM[252] =	32'b00000000000000000000000000111111;
    RAM[253] =	32'b00000000000000000000000000111111;
    RAM[254] =	32'b00000000000000000000000000111111;
    RAM[255] =	32'b00000000000000000000000000111111;
    RAM[256] =	32'b00000000000000000000000000111111;
    RAM[257] =	32'b00000000000000000000000000111111;
    RAM[258] =	32'b00000000000000000000000000111111;
    RAM[259] =	32'b00000000000000000000000000111111;
    RAM[260] =	32'b00000000000000000000000000111111;
    RAM[261] =	32'b00000000000000000000000000111111;
    RAM[262] =	32'b00000000000000000000000000111111;
    RAM[263] =	32'b00000000000000000000000000010000;
    RAM[264] =	32'b00000000000000000000000000010000;
    RAM[265] =	32'b00000000000000000000000000111111;
    RAM[266] =	32'b00000000000000000000000000111111;
    RAM[267] =	32'b00000000000000000000000000111111;
    RAM[268] =	32'b00000000000000000000000000111111;
    RAM[269] =	32'b00000000000000000000000000111111;
    RAM[270] =	32'b00000000000000000000000000111111;
    RAM[271] =	32'b00000000000000000000000000111111;
    RAM[272] =	32'b00000000000000000000000000111111;
    RAM[273] =	32'b00000000000000000000000000111111;
    RAM[274] =	32'b00000000000000000000000000111111;
    RAM[275] =	32'b00000000000000000000000000111111;
    RAM[276] =	32'b00000000000000000000000000111111;
    RAM[277] =	32'b00000000000000000000000000111111;
    RAM[278] =	32'b00000000000000000000000000111111;
    RAM[279] =	32'b00000000000000000000000000111111;
    RAM[280] =	32'b00000000000000000000000000111111;
    RAM[281] =	32'b00000000000000000000000000111111;
    RAM[282] =	32'b00000000000000000000000000111111;
    RAM[283] =	32'b00000000000000000000000000111111;
    RAM[284] =	32'b00000000000000000000000000111111;
    RAM[285] =	32'b00000000000000000000000000111111;
    RAM[286] =	32'b00000000000000000000000000111111;
    RAM[287] =	32'b00000000000000000000000000111111;
    RAM[288] =	32'b00000000000000000000000000111111;
    RAM[289] =	32'b00000000000000000000000000111111;
    RAM[290] =	32'b00000000000000000000000000111111;
    RAM[291] =	32'b00000000000000000000000000111111;
    RAM[292] =	32'b00000000000000000000000000111111;
    RAM[293] =	32'b00000000000000000000000000111111;
    RAM[294] =	32'b00000000000000000000000000000011;
    RAM[295] =	32'b00000000000000000000000000001100;
    RAM[296] =	32'b00000000000000000000000000110000;
    RAM[297] =	32'b00000000000000000000000000111100;
    RAM[298] =	32'b00000000000000000000000000110011;
    RAM[299] =	32'b00000000000000000000000000001111;
  end

  assign vdata = RAM[vaddr[31:0]]; 
  assign read_data = RAM[addr[31:2]]; // word aligned
  
  always_ff @(posedge clk) 
    if (mem_write) 
	 begin
		RAM[addr[31:2]] 		<= write_data;
	end
endmodule

// Modulo de memoria das instruçoes
module imem(input  logic [31:0] pc,
            output logic [31:0] instr);

  logic [31:0] RAM[32:0];
 
  initial begin
		RAM[0]  = 32'h00000493;
		RAM[1]  = 32'h0200006f;
		RAM[2]  = 32'h000007b7;
		RAM[3]  = 32'h00078713;
		RAM[4]  = 32'h00249793;
		RAM[5]  = 32'h00f707b3;
		RAM[6]  = 32'h00f00713;
		RAM[7]  = 32'h00e7a023;
		RAM[8]  = 32'h00148493;
		RAM[9]  = 32'h000027b7;
		RAM[10] = 32'h00078793;
		RAM[11] = 32'h57f78793;
		RAM[12] = 32'hfc97dce3;
		RAM[13] = 32'h00000793;
		RAM[14] = 32'h00f00533;
		RAM[15] = 32'h00008067;
  end
  

  assign instr = RAM[pc[31:2]]; // word aligned
endmodule